module tx_baud_rate_generator(
    input tx_clk,
    input [1:0] tx_sel,
    output reg tx_baud_out;
);

    wire 
endmodule

`ifndef UART_PARAMS

`define UART_PARAMS

`ifndef DATA_WIDTH 
    `define DATA_WIDTH 8
`endif
`endif
